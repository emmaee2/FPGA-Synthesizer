//module fir_filter(
//		input [(LN):0] sample,
//		output [(LN):0] average
//)
//parameter LN = 16;
//
//
//
//endmodule
